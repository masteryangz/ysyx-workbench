module led(
  input clk,
  input rst,
  input [4:0] btn,
  input [15:0] sw,
  output [2:0] ledr
);

//  assign ledr[0] = ready;
//  assign ledr[1] = sampling;
//  assign ledr[2] = overflow;

endmodule
